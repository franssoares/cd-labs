library verilog;
use verilog.vl_types.all;
entity ffd_6_vlg_vec_tst is
end ffd_6_vlg_vec_tst;
