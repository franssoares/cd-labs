library verilog;
use verilog.vl_types.all;
entity reg_8x1_vlg_vec_tst is
end reg_8x1_vlg_vec_tst;
