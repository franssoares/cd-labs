library verilog;
use verilog.vl_types.all;
entity RF_16x16_vlg_vec_tst is
end RF_16x16_vlg_vec_tst;
