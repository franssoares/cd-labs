library verilog;
use verilog.vl_types.all;
entity FFD_vlg_vec_tst is
end FFD_vlg_vec_tst;
