library verilog;
use verilog.vl_types.all;
entity divide_freq_vlg_vec_tst is
end divide_freq_vlg_vec_tst;
