library verilog;
use verilog.vl_types.all;
entity ffd_5_vlg_vec_tst is
end ffd_5_vlg_vec_tst;
