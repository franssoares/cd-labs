library verilog;
use verilog.vl_types.all;
entity bf_8x1_vlg_vec_tst is
end bf_8x1_vlg_vec_tst;
