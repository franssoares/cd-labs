library verilog;
use verilog.vl_types.all;
entity datapath_control_vlg_vec_tst is
end datapath_control_vlg_vec_tst;
