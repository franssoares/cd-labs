library verilog;
use verilog.vl_types.all;
entity reg_1x5_vlg_vec_tst is
end reg_1x5_vlg_vec_tst;
