library verilog;
use verilog.vl_types.all;
entity counter_wload_6_vlg_vec_tst is
end counter_wload_6_vlg_vec_tst;
