library verilog;
use verilog.vl_types.all;
entity unid_control_vlg_vec_tst is
end unid_control_vlg_vec_tst;
