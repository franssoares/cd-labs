library verilog;
use verilog.vl_types.all;
entity calculadora_vlg_vec_tst is
end calculadora_vlg_vec_tst;
