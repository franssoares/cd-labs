library verilog;
use verilog.vl_types.all;
entity timer_vlg_vec_tst is
end timer_vlg_vec_tst;
