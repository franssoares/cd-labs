library verilog;
use verilog.vl_types.all;
entity controle_vlg_vec_tst is
end controle_vlg_vec_tst;
