library verilog;
use verilog.vl_types.all;
entity controlador_vlg_vec_tst is
end controlador_vlg_vec_tst;
