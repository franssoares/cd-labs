library verilog;
use verilog.vl_types.all;
entity counter_min_6_vlg_vec_tst is
end counter_min_6_vlg_vec_tst;
