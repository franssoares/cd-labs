library verilog;
use verilog.vl_types.all;
entity ula_vlg_vec_tst is
end ula_vlg_vec_tst;
