library verilog;
use verilog.vl_types.all;
entity counter_seg_6_vlg_vec_tst is
end counter_seg_6_vlg_vec_tst;
