library verilog;
use verilog.vl_types.all;
entity LatchD_vlg_vec_tst is
end LatchD_vlg_vec_tst;
