-- Biblioteca
LIBRARY ieee;
USE ieee.std_logic_1164.all;
	 
-- Entidade
ENTITY bf_8x22 is
    port (
		w_data : in std_logic_vector(21 downto 0);
		w_addr : in STD_LOGIC_VECTOR(2 DOWNTO 0);
		w_en : in std_logic;
		r_data : out std_logic_vector(21 downto 0);
		r_addr : in STD_LOGIC_VECTOR(2 DOWNTO 0);
		r_en : in std_logic;
		
	    clk : in std_logic;
		en :  in std_logic;              
		clear : in std_logic;						
		load : in std_logic
	);
END ENTITY bf_8x22;

-- Arquitetura
ARCHITECTURE behav OF bf_8x22 IS

-- Componentes

	-- Registrador
	COMPONENT reg_8x22 is
		port (
			d_data : in std_logic_vector(21 downto 0);        -- Entrada de dados
			clk : in std_logic;                 -- Sinal de clock
			clear : in std_logic;						-- Sinal de clear
			load : in std_logic; 		  				-- Sinal de carga
			q_data : out std_logic_vector(21 downto 0)
		);
	END COMPONENT reg_8x22;

	--Decoder
	COMPONENT dcd_3x8 is
		PORT(
			in_id : STD_LOGIC_VECTOR(2 DOWNTO 0); -- ID
        	en : STD_LOGIC; --ENABLE
			d : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT dcd_3x8;

	-- Driver de 3 estados
	COMPONENT tri_states_driver_22 IS
		PORT(
			in_data : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
			enable : IN STD_LOGIC;
			out_data : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
		);
	END COMPONENT tri_states_driver_22;

-- Fios

	SIGNAL decoder0_wires : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL decoder1_wires : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL reg0_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg1_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg2_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg3_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg4_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg5_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg6_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	SIGNAL reg7_wires : STD_LOGIC_VECTOR(21 DOWNTO 0);
	
BEGIN

    -- Instancia
    decoder1 : dcd_3x8
    PORT MAP(
      in_id => w_addr,
	   en => w_en,
	   d => decoder0_wires
    );

	reg0_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(0),
		q_data => reg0_wires
	);
	
	reg1_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(1),
		q_data => reg1_wires
	);
	
	reg2_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(2),
		q_data => reg2_wires
	);
	
	reg3_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(3),
		q_data => reg3_wires
	);
	
	reg4_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(4),
		q_data => reg4_wires
	);
	
	reg5_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(5),
		q_data => reg5_wires
	);
	
	reg6_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(6),
		q_data => reg6_wires
	);
	
	reg7_1x22 : reg_8x22
	PORT MAP(
		d_data => w_data,
		clk => clk,
		clear => clear,
		load => decoder0_wires(7),
		q_data => reg7_wires
	);

	tsd0 : tri_states_driver_22
	PORT MAP(
		in_data => reg0_wires,
		enable => decoder1_wires(0),
		out_data => r_data
	);
	
	tsd1 : tri_states_driver_22
	PORT MAP(
		in_data => reg1_wires,
		enable => decoder1_wires(1),
		out_data => r_data
	);
	
	tsd2 : tri_states_driver_22
	PORT MAP(
		in_data => reg2_wires,
		enable => decoder1_wires(2),
		out_data => r_data
	);
	
	tsd3 : tri_states_driver_22
	PORT MAP(
		in_data => reg3_wires,
		enable => decoder1_wires(3),
		out_data => r_data
	);
	
	tsd4 : tri_states_driver_22
	PORT MAP(
		in_data => reg4_wires,
		enable => decoder1_wires(4),
		out_data => r_data
	);
	
	tsd5 : tri_states_driver_22
	PORT MAP(
		in_data => reg5_wires,
		enable => decoder1_wires(5),
		out_data => r_data
	);
	
	tsd6 : tri_states_driver_22
	PORT MAP(
		in_data => reg6_wires,
		enable => decoder1_wires(6),
		out_data => r_data
	);
	
	tsd7 : tri_states_driver_22
	PORT MAP(
		in_data => reg7_wires,
		enable => decoder1_wires(7),
		out_data => r_data
	);
	
	decoder2 : dcd_3x8
	PORT MAP(
		in_id => r_addr,
		en => r_en,
		d => decoder1_wires
	);

END ARCHITECTURE behav;