library verilog;
use verilog.vl_types.all;
entity reg_1x6_vlg_vec_tst is
end reg_1x6_vlg_vec_tst;
