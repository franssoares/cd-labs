library verilog;
use verilog.vl_types.all;
entity bf_8x22_vlg_vec_tst is
end bf_8x22_vlg_vec_tst;
