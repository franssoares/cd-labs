library verilog;
use verilog.vl_types.all;
entity datapath_vlg_vec_tst is
end datapath_vlg_vec_tst;
