library verilog;
use verilog.vl_types.all;
entity comb_logic_vlg_vec_tst is
end comb_logic_vlg_vec_tst;
